*** SPICE deck for cell not{lay} from library Digital
*** Created on Sat Apr 24, 2021 12:22:30
*** Last revised on Sat Apr 24, 2021 12:45:41
*** Written on Sat Apr 24, 2021 12:46:07 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*** WARNING: no ground connection for N-transistor wells in cell 'not{lay}'

*** TOP LEVEL CELL: not{lay}
Mnmos@0 vss vin vout gnd NMOS L=0.6U W=3U AS=8.1P AD=9.9P PS=12.6U PD=18.6U
Mpmos@0 vdd vin vout vss PMOS L=0.6U W=6U AS=8.1P AD=19.8P PS=12.6U PD=30.6U

* Spice Code nodes in cell cell 'not{lay}'
.include D:\Electric\C5_models.txt
vdd vdd 0 DC 5
vss vss 0 DC 0
vin vin 0 pulse(0 5 0 1n 1n 10n 20n)
.trans 0 40n
.END
