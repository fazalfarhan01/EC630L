*** SPICE deck for cell nor{lay} from library Digital
*** Created on Sat Apr 24, 2021 14:15:00
*** Last revised on Sat Apr 24, 2021 14:27:17
*** Written on Sat Apr 24, 2021 14:27:34 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*** WARNING: no ground connection for N-transistor wells in cell 'nor{lay}'

*** TOP LEVEL CELL: nor{lay}
Mnmos@0 vss vin1 vout gnd NMOS L=0.6U W=3U AS=7.2P AD=7.65P PS=11.6U PD=14.1U
Mnmos@1 vout vin2 vss gnd NMOS L=0.6U W=3U AS=7.65P AD=7.2P PS=14.1U PD=11.6U
Mpmos@0 net@1 vin1 vdd vss PMOS L=0.6U W=6U AS=19.8P AD=10.8P PS=30.6U PD=15.6U
Mpmos@1 vout vin2 net@1 vss PMOS L=0.6U W=6U AS=10.8P AD=7.2P PS=15.6U PD=11.6U

* Spice Code nodes in cell cell 'nor{lay}'
.include D:\Electric\C5_models.txt 
vdd vdd 0 DC 5
vss vss 0 DC 0
vin1 vin1 0 pulse 5 0 0 1n 1n 2u 4u
vin2 vin2 0 pulse 5 0 0 1n 1n 1u 2u
.tran 4u
.END
