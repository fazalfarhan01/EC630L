*** SPICE deck for cell nand{lay} from library Digital
*** Created on Sat Apr 24, 2021 13:26:23
*** Last revised on Sat Apr 24, 2021 14:01:29
*** Written on Sat Apr 24, 2021 14:01:43 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*** WARNING: no ground connection for N-transistor wells in cell 'nand{lay}'

*** TOP LEVEL CELL: nand{lay}
Mnmos@0 net@3 vin1 vout gnd NMOS L=0.6U W=3U AS=9P AD=5.4P PS=13.6U PD=9.6U
Mnmos@1 vss vin2 net@3 gnd NMOS L=0.6U W=3U AS=5.4P AD=10.8P PS=9.6U PD=19.2U
Mpmos@0 vdd vin1 vout vss PMOS L=0.6U W=6U AS=9P AD=15.3P PS=13.6U PD=23.1U
Mpmos@1 vout vin2 vdd vss PMOS L=0.6U W=6U AS=15.3P AD=9P PS=23.1U PD=13.6U

* Spice Code nodes in cell cell 'nand{lay}'
.include D:\Electric\C5_models.txt 
vdd vdd 0 DC 5
vss vss 0 DC 0
vin1 vin1 0 pulse 5 0 0 1n 1n 2u 4u
vin2 vin2 0 pulse 5 0 0 1n 1n 1u 2u
.tran 4u
.END
