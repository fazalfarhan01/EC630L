*** SPICE deck for cell NAND{lay} from library NAND
*** Created on Fri Apr 23, 2021 15:47:53
*** Last revised on Fri Apr 23, 2021 22:16:22
*** Written on Fri Apr 23, 2021 22:16:34 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: NAND{lay}
Mnmos@0 net@4 A vout vss NMOS L=0.6U W=3U AS=8.25P AD=4.95P PS=13.3U PD=9.3U
Mnmos@1 vss B net@4 vss NMOS L=0.6U W=3U AS=4.95P AD=9.45P PS=9.3U PD=18.3U
Mpmos@0 vdd A vout vdd PMOS L=0.6U W=6U AS=8.25P AD=14.4P PS=13.3U PD=22.8U
Mpmos@1 vdd B vout vdd PMOS L=0.6U W=6U AS=8.25P AD=14.4P PS=13.3U PD=22.8U

* Spice Code nodes in cell cell 'NAND{lay}'
.include D:\Electric\C5_models.txt 
vdd vdd 0 DC 5
vss vss 0 DC 0
Va A 0 pulse 5 0 0 1n 1n 2u 4u
Vb B 0 pulse 5 0 0 1n 1n 1u 2u
.tran 4u
.END
